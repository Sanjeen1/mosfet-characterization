.include ./tsmc180.txt

m1 vdd in 0 0 nfet w=3u l=0.5u
v_dd vdd 0 3.3
v_in in 0 3.3
.dc v_dd 0 3.3 0.1 v_in 0 3.3 1
.control
foreach lam .01 .1 10
altermod m1 PCLM = $lam
run

end
.endc
.control
foreach iter 1 2 3

setplot dc$iter
plot -v_dd#branch
end

set color0=white
set color1=black
set color2=red

set xbrushwidth=3
.endc
.end