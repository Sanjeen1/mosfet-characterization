.include ./t14y.txt
.Temp 27

m1 vdd in 0 0 CMOSN w=10u l=3u
v_dd vdd 0 3.3
v_in in 0 3.3

.dc v_in 0 3.3 0.1
.control
foreach t 20 50 100
alter m1 Temp = $t
run
end
.endc
.control
foreach iter 1 2 3
setplot dc$iter
plot -v_dd#branch 
end
set color0=white
set color1=black
set color2=red
set color2=pink
set xbrushwidth=3

plot dc1.v_dd#branch*-1 dc2.v_dd#branch*-1 dc3.v_dd#branch*-1
.endc

.end