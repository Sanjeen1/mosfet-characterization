.include ./tsmc180.txt
m1 vdd in 0 0 nfet w=10u l=3u
v_dd vdd 0 3.3
v_in in 0 3.3
.dc v_in 0 3.3 0.1 v_dd 0 2 2

.control
foreach vt 0.1 0.4 
altermod m1 VTH0 = $vt
run
end
.endc
.control
foreach iter 1 2 

setplot dc$iter
plot -v_dd#branch 
end
set color0=white
set color1=black
set color2=red

set xbrushwidth=3
  print v(vdd)
 

.endc
.end