.include ./tsmc180.txt

m1 vdd in s 0 nfet w=10u l=3u
v_dd vdd 0 3.3
v_in in 0 3.3

v_sb s 0 1.8

.dc v_in 0 3.3 0.1 v_sb 0 1.8 0.6
.control
run

plot -v_dd#branch

set color0=white
set color1=black
set color2=blue

set xbrushwidth=3
.endc
.end