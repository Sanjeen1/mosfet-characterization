.include ./tsmc180.txt

m1 vdd in 0 0 nfet w=3u l=3u

v_dd vdd 0 5
v_in in 0 5
.dc v_dd 0 5 0.1 v_in 0 5 1

.control
foreach dim 0.1u 5u 10u
alter m1 w = $dim
run
end
.endc
.control
foreach iter 1 2 3

setplot dc$iter
plot -v_dd#branch

end

set color0=white
set color1=black
set color2=red

set xbrushwidth=3

.endc
.end